* C:\Users\Acer\eSim-Workspace\abdulmannan\abdulmannan.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/04/22 11:56:32

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  io i1 set Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ adc_bridge_3		
U6  Net-_U4-Pad4_ Net-_SC1-Pad1_ dac_bridge_1		
v3  set GND pulse		
v2  i1 GND pulse		
v1  io GND pulse		
U3  set plot_db		
U2  i1 plot_db		
U1  io plot_db		
SC2  vout GND sky130_fd_pr__cap_mim_m3_1		
U7  vout plot_db		
scmode1  SKY130mode		
SC1  Net-_SC1-Pad1_ vout Net-_SC1-Pad1_ sky130_fd_pr__res_generic_pd		
U8  ? ? ? ? abdulmannan_mux		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ abdulmannan_mux		

.end
